module regfile(
	input 
	);



endmodule
