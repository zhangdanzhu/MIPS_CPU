~timescale 1ns / 1ps

module pipeline_mips_cpu(
	input clk
	output xxx
	);

	wire 


endmodule
